module led(F, D);
input [3:0] D;
output [6:0]F;
reg [6:0]F;
//wire [6:0]F;


always@(D)
case(D)
4'b0000:F<=7'b1000000;//0
4'b0001:F<=7'b1111001;//1
4'b0010:F<=7'b0100100;//2
4'b0011:F<=7'b0110000;//3
4'b0100:F<=7'b0011001;//4
4'b0101:F<=7'b0010010;//5
4'b0110:F<=7'b0000010;//6
4'b0111:F<=7'b1111000;//7
4'b1000:F<=7'b0000000;//8
4'b1001:F<=7'b0010000;//9
    default: F<=7'b1111111;
endcase
endmodule

 