module tb_74LS138; 
    wire [6:0]F; 
    reg [3:0]D;
   led   dec(F,D);
initial begin
$monitor("%b,%b,%b,%b,%b,%b,%b",F[0],F[1],F[2],F[3],F[4],F[5],F[6]); 
$display("%3t: D0 = %b, D1 = %b, D2=%b, D3=%b, F1=%b, F2=%b, F3=%b, F4=%b, F5 = %b, F6=%b, F7=%b",$time,D[0],D[1],D[2],D[3],F[0],F[1],F[2],F[3],F[4],F[5],F[6]); 
 #5 D[0]=0; D[1]=0; D[2]=0; D[3]=0;//0
 #5 D[0]=1; D[1]=0; D[2]=0; D[3]=0;//1
 #5 D[0]=0; D[1]=1; D[2]=0; D[3]=0;//2
 #5 D[0]=1; D[1]=1; D[2]=0; D[3]=0;//3
 #5 D[0]=0; D[1]=0; D[2]=1; D[3]=0;//4
 #5 D[0]=1; D[1]=0; D[2]=1; D[3]=0;//5
 #5 D[0]=0; D[1]=1; D[2]=1; D[3]=0;//6
 #5 D[0]=1; D[1]=1; D[2]=1; D[3]=0;//7
 #5 D[0]=0; D[1]=0; D[2]=0; D[3]=1;//8
 #5 D[0]=1; D[1]=0; D[2]=0; D[3]=1;//9
 #5 D[0]=1; D[1]=0; D[2]=1; D[3]=1;//其他

 
  #10 $finish; 
  end 
   endmodule