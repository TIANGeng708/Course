module kmap(F, A, B, C, D);
input A, B, C, D;
output F;
wire notA, notB, notC, notD;
wire and1, and2, and3;
//F=B'D'+CD'+ABC'D
not not_1 (notA, A);
not not_1 (notB, B);
not not_1 (notC, C);
not not_1 (notD, D);
and and_1 (anda, C, notD);
and and_2 (andb, notB, notD);
and and_3 (andc, A, B, notC, D);
or or_1 (F, anda, andb, andc);


endmodule
module kmap1;
reg a, b, c, d;
wire f;

kmap com_1(f, a, b, c, d);

initial begin
 $monitor("%3t: a is %b, b is %b, c is %b, d %b, f is %b.", $time, a, b, c, d, f);
  # 5 a = 1; b = 0; c=0; d=0;
  # 5 a = 1; b = 1; c=0; d=0;
  # 5 a = 1; b = 0; c=1; d=0;
  # 5 a = 1; b = 0; c=0; d=1;
  # 5 a = 1; b = 1; c=1; d=0;
  # 5 a = 1; b = 1; c=0; d=1;
  # 5 a = 1; b = 0; c=1; d=1;
  # 5 a = 1; b = 1; c=1; d=1;
  # 5 a = 0; b = 0; c=0; d=0;
  # 5 a = 0; b = 1; c=0; d=0;
  # 5 a = 0; b = 0; c=1; d=0;
  # 5 a = 0; b = 0; c=0; d=1;
  # 5 a = 0; b = 1; c=1; d=0;
  # 5 a = 0; b = 1; c=0; d=1;
  # 5 a = 0; b = 0; c=1; d=1;
  # 5 a = 0; b = 1; c=1; d=1;
  # 10 $finish; 
 end 
 endmodule