module test_tb; 

wire [31:0]Q;
wire  [31:0]R;
reg [31:0]A;
reg [31:0]B;
reg CLK;
reg reset;


divide myadd(Q, R, A, B,CLK,reset);
initial begin
    A=32'b01110010000000000000000000000000;
end
initial begin
    B=32'b00000000000000000000000000000100;
end
initial begin
    CLK=1'b1;
end
initial begin
    reset=1'b1;
end
always@(CLK)
begin
    #1 CLK<=!CLK;
end

always@(reset)
begin
    #3 reset<=!reset;
end

initial begin 
$monitor("%3t:%b   %b   %b   %b ",$time,A,B,Q,R,CLK,reset); 
# 3 A=32'b00000010000000000000000000000000;B=32'b00000000000000000000000000000100;
# 3 A=32'b00000010000000000000000000000000;B=32'b00000000000000000000000000000010;
# 3 A=32'b00000010000000000000000000000000;B=32'b00000000000000000000000000100000;
# 3 A=32'b00000010000000000000011100000000;B=32'b00000000000000000000000000000110;
# 3 A=32'b00110010000000000000000000000100;B=32'b00000000000000000011111110000010;
# 3 A=32'b00000011010000000000011100000000;B=32'b00000000000000000000011100100000;
# 100 $finish;
  end 
  endmodule